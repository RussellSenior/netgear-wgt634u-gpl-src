Template: ifupdown/convert-interfaces
Type: boolean
Default: true
Description: Update /etc/network/interfaces?
 The format of /etc/network/interfaces has had a minor but incompatible
 change made between version 0.5.x and 0.6.x of ifupdown. It is however
 possible to automatically convert from the old format to the new in almost
 all cases.
Description-sv: Uppdatera /etc/network/interfaces?
 Formatet p� /etc/network/interfaces genomgick en liten men inkompatibel
 �ndring mellan version 0.5.x och 0.6.x av ifupdown. Det �r dock m�jligt
 att n�stan alltid automatiskt konvertera fr�n det gamla formatet
 till det nya.
